.Addotional power values for 3D IC Thermal Grid (3x3x3 = 27 nodes)

.--- Fixed temperature sources ---
VAMB3 0_2_0 0 300
VAMB4 2_0_2 0 300

.--- Power sources ---
I7 0 2_2_2 1

.print dc v(*)
.op
.end