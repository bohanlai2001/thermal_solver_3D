.3D IC Thermal Grid (3x3x3 = 27 nodes)
.Node naming: X_Y_Z (0-based indices)
.Resistors numbered sequentially (R1, R2, ...)

.--- Resistances (adjacent nodes connected) ---
R1  0_0_0 1_0_0 1
R2  1_0_0 2_0_0 1
R3  0_1_0 1_1_0 1
R4  1_1_0 2_1_0 1
R5  0_2_0 1_2_0 1
R6  1_2_0 2_2_0 1
R7  0_0_1 1_0_1 1
R8  1_0_1 2_0_1 1
R9  0_1_1 1_1_1 1
R10 1_1_1 2_1_1 1
R11 0_2_1 1_2_1 1
R12 1_2_1 2_2_1 1
R13 0_0_2 1_0_2 1
R14 1_0_2 2_0_2 1
R15 0_1_2 1_1_2 1
R16 1_1_2 2_1_2 1
R17 0_2_2 1_2_2 1
R18 1_2_2 2_2_2 1
R19 0_0_0 0_1_0 1
R20 0_1_0 0_2_0 1
R21 1_0_0 1_1_0 1
R22 1_1_0 1_2_0 1
R23 2_0_0 2_1_0 1
R24 2_1_0 2_2_0 1
R25 0_0_1 0_1_1 1
R26 0_1_1 0_2_1 1
R27 1_0_1 1_1_1 1
R28 1_1_1 1_2_1 1
R29 2_0_1 2_1_1 1
R30 2_1_1 2_2_1 1
R31 0_0_2 0_1_2 1
R32 0_1_2 0_2_2 1
R33 1_0_2 1_1_2 1
R34 1_1_2 1_2_2 1
R35 2_0_2 2_1_2 1
R36 2_1_2 2_2_2 1
R37 0_0_0 0_0_1 1
R38 0_0_1 0_0_2 1
R39 1_0_0 1_0_1 1
R40 1_0_1 1_0_2 1
R41 2_0_0 2_0_1 1
R42 2_0_1 2_0_2 1
R43 0_1_0 0_1_1 1
R44 0_1_1 0_1_2 1
R45 1_1_0 1_1_1 1
R46 1_1_1 1_1_2 1
R47 2_1_0 2_1_1 1
R48 2_1_1 2_1_2 1
R49 0_2_0 0_2_1 1
R50 0_2_1 0_2_2 1
R51 1_2_0 1_2_1 1
R52 1_2_1 1_2_2 1
R53 2_2_0 2_2_1 1
R54 2_2_1 2_2_2 1

.--- Fixed temperature sources ---
VAMB1 0_0_0 0 300
VAMB2 2_2_2 0 300

.--- Power sources ---
I1 0 1_1_0 1
I2 0 0_2_1 1
I3 0 1_0_2 1
I4 0 2_1_1 1
I5 0 1_2_2 1
I6 0 2_0_2 1

.print dc v(*)
.op
.end